

// `ifndef __CHECKER_COMMON__
// `define __CHECHER_COMMON__

// `include "uart_uvc.svh"

// class checkr_comm;
// 	static int unsigned err_cnt;
// endclass : checkr_comm

// `endif // __CHECKER_COMMON__

// `ifndef __UART_TRANSMIT_CHECKER__
// `define __UART_TRANSMIT_CHECKER__

// class uart_check;
	
// endclass : uart_check

// `endif //__UART_TRANSMIT_CHECKER__