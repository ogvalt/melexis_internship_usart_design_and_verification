module transmitter	(
					i_txclk,
					i_rst_n,	
					i_tx_data,
					i_tx_data_9bit,
					i_tx_data_en,
					i_ucz,
					i_upm,
					i_usbs,
					o_tx,
					o_transmit_complete,
					o_data_read_from_udr
					);

/*--------------------------Parameter--------------------------*/

/*--------------------------Input ports------------------------*/

input 					i_txclk; 		// clock signal for transmitter1 ggenerated by Clock Generator
input 					i_rst_n;		// system reset

input 	[7:0]			i_tx_data;		// data from UDR(transmit)
input 					i_tx_data_9bit;	// 9th bit for transmitter1
input 					i_tx_data_en; 	// new data for transmit enable, 

input 	[2:0]			i_ucz;			// character size 
	/*	
		|UCZ2	|UCZ1	|UCZ0	|Character size		|
	 	|	0	|	0	|	0	|	5-bit			|
	 	|	0	|	0	|	1	|	6-bit			|
	 	|	0	|	1	|	0	|	7-bit			|
	 	|	0	|	1	|	1	|	8-bit			|
	 	|	1	|	0	|	0	|	Reserved		|
	 	|	1	|	0	|	1	|	Reserved		|
	 	|	1	|	1	|	0	|	Reserved		|
	 	|	1	|	1	|	1	|	9-bit			|
	*/

input 	[1:0]			i_upm;			//	parity mode
	/*
		|UPM1	|UPM0	|Parity mode 	|
		|	0	|	0	|Disable		|
		|	0	|	1	|Reserved		|
		|	1	|	0	|Enable, Even	|
		|	1	|	1	|Enable, Odd	|
	*/

input 					i_usbs; 		// stop bit select, 0 - 1-bit, 1 - 2-bit

/*--------------------------Ouput ports------------------------*/

output					o_transmit_complete;	// transmit complete flag
												// it will use as empty flag, that will overwrite
												// UDR empty flag
output  reg 			o_tx;					// tx line
output 					o_data_read_from_udr;

/*--------------------------Inout ports------------------------*/

/*--------------------------Variables--------------------------*/

reg		[8:0]			shift_register; // transmit shift register

reg 	[3:0]			counter;

wire 					fsm_start_bit; 		  // start bit insert signal

wire					fsm_rewrite_or_shift; // rewrite or shift transmit shift register
										  	  // 1-rewrite, 0 - shift
wire 					fsm_counter_en;		  // 1 - counter rewrite, 0 - counting
wire					fsm_parity_generate;  // signal to parity checker to generate parity bit
wire 					fsm_parity_insert;	  // signal that enables parity insert
wire 					fsm_stop_bit_insert;  // stop bit signal insert
wire 					fsm_transmit_complete;// transmit complete
wire  					fsm_data_transmit;	  // data in transmit process signal

wire 					last_bit_flag;			  // counter = 0, so last bit is sent

wire					parity_bit;			  // parity bit gets from parity checker

reg 					parity_bit_reg; 	  

wire 					tx;
reg 					data_read_from_udr;

/*--------------------------Modules Instances-------------------*/

parity_checker  parity_check1 (
				              	.i_clk 				(i_txclk),
				              	.i_rst_n			(i_rst_n),  
				              	.i_parity_mode_0	(i_upm[0]),
				              	.i_parity_en		(fsm_parity_generate),
				              	.i_frame_size		(i_ucz),
				              	.i_frame 			({i_tx_data_9bit, i_tx_data}),
				              	.o_parity_check		(parity_bit)
				              );

fsm_tx 	transmitter1_fsm1	( 
								.i_txclk				(i_txclk), 
								.i_rst_n				(i_rst_n),
								.i_data_in_udr			(i_tx_data_en),
								.i_last_bit_sent		(last_bit_flag),
								.i_upm1					(i_upm[1]),
								.i_usbs					(i_usbs),
								.o_start_bit_insert		(fsm_start_bit),
								.o_parity_generate		(fsm_parity_generate),
				    			.o_reg_wr_or_shift		(fsm_rewrite_or_shift),
				    			.o_rewr_or_count		(fsm_counter_en),
				    			.o_data_transmit		(fsm_data_transmit),
				    			.o_parity_insert		(fsm_parity_insert),
				    			.o_stop_bit				(fsm_stop_bit_insert),
				    			.o_transmit_complete	(fsm_transmit_complete)
				              );

/*--------------------------Sequential logic-------------------*/
assign  o_data_read_from_udr = data_read_from_udr;
assign 	last_bit_flag	=	(counter == 1);
assign 	o_transmit_complete = fsm_transmit_complete;
assign  tx 				= shift_register[0];

/*--------------------------Combinational logic----------------*/


always @(posedge i_txclk or negedge i_rst_n) begin : shift_register_load_block
	if(~i_rst_n) begin : shift_register_reset
		shift_register <= 0;
		data_read_from_udr <= 0;
	end else begin : shift_register_operation
		if (fsm_rewrite_or_shift) begin	
			shift_register <= {i_tx_data_9bit, i_tx_data};
			data_read_from_udr <= 1;
		end else begin
			data_read_from_udr <= 0;
			shift_register <= {1'b0, shift_register[8:1]};
		end
	end
end // shift_register_load_block

always @(posedge i_txclk or negedge i_rst_n) begin : proc_
	if(~i_rst_n) begin
		parity_bit_reg <= 0;
	end else begin
		if (fsm_parity_generate) 
			parity_bit_reg <= parity_bit;
	end
end

always @(posedge i_txclk or negedge i_rst_n) begin : counter_block
	if(~i_rst_n) begin : counter_reset
		counter <= 0;
	end else begin : counter_operation
		if (fsm_counter_en|!fsm_data_transmit) begin
			case(i_ucz)
				3'b000:		counter <= 5; // 5-bit  
				3'b001:		counter <= 6; // 6-bit
				3'b010:		counter <= 7; // 7-bit
				3'b011:		counter <= 8; // 8-bit
				3'b111:		counter <= 9; // 9-bit
				default:	counter <= 0; // Reserved
			endcase // i_ucz
		end else begin
			counter <= counter - 1;
		end
	end
end

always @(posedge i_txclk or negedge i_rst_n) begin : tx_line_block
	if(~i_rst_n) begin
		o_tx <= 1;
	end else begin
		if (fsm_parity_insert)	o_tx <= parity_bit_reg;
		else begin
			if (fsm_stop_bit_insert) 		o_tx <= 1;
			else begin
				if (fsm_start_bit) 			o_tx <= 0;
				else begin
					if (fsm_data_transmit) 	o_tx <= tx;
					else 					o_tx <= 1;
				end
			end
		end
	end
end // tx_line_block



/*--------------------------Finite state machine---------------*/

endmodule